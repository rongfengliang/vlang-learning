
module main

import fetchbaidu

fn main() {

    fetchbaidu.fetchindexpage()
}